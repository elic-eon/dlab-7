//Subject:
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      Szuyi Huang
//----------------------------------------------
//Date:        2013-12-11 13:39
//----------------------------------------------
//Description:
//--------------------------------------------------------------------------------
module radius_control(

					);

//--------------------------------------------------------------------------------
// I/O ports declearation


//--------------------------------------------------------------------------------
// Internal signal

//--------------------------------------------------------------------------------
// Parameter declearation

endmodule

